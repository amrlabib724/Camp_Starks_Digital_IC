
module And2 (A,B,C);
  input A,B;
  output C;
  assign y=A&B;
    
endmodule